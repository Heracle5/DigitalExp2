module counter(
    
);

endmodule