module LogicProcessingUnited();

endmodule